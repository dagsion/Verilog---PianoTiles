module audio (
	// Inputs
	CLOCK_50,
	KEY,

	AUD_ADCDAT,

	// Bidirectionals
	AUD_BCLK,
	AUD_ADCLRCK,
	AUD_DACLRCK,

	FPGA_I2C_SDAT,

	// Outputs
	AUD_XCK,
	AUD_DACDAT,

	FPGA_I2C_SCLK,
	SW,
	
	PS2_CLK,					// PS2 Clock
	PS2_DAT
);

/*****************************************************************************
 *                           Parameter Declarations                          *
 *****************************************************************************/


/*****************************************************************************
 *                             Port Declarations                             *
 *****************************************************************************/
// Inputs
input				CLOCK_50;
input				[3:0]KEY;
input 			[3:0]SW;

input				AUD_ADCDAT;

// Bidirectionals
inout				AUD_BCLK;
inout				AUD_ADCLRCK;
inout				AUD_DACLRCK;

inout				FPGA_I2C_SDAT;

inout 			PS2_CLK;					// PS2 Clock
inout				PS2_DAT;

// Outputs
output				AUD_XCK;
output				AUD_DACDAT;

output				FPGA_I2C_SCLK;



/*****************************************************************************
 *                 Internal Wires and Registers Declarations                 *
 *****************************************************************************/
// Internal Wires
wire				audio_in_available;
wire		[31:0]	left_channel_audio_in;
wire		[31:0]	right_channel_audio_in;
wire				read_audio_in;

wire				audio_out_allowed;
wire		[31:0]	left_channel_audio_out;
wire		[31:0]	right_channel_audio_out;
wire				write_audio_out;

wire 		[7:0]keyboard;
wire 		e;

// Internal Registers

reg [18:0] delay_cnt;
reg [18:0] delay;

reg snd;

// State Machine Registers

/*****************************************************************************
 *                         Finite State Machine(s)                           *
 *****************************************************************************/
 
always @(posedge e)
begin
	case(keyboard)
	8'b00010101: delay<=32'h2F691;
	8'b00011101: delay<=32'h29AB2;
	8'b00100100: delay<=32'h24A26;
	8'b00101101: delay<=32'h230E4;
	8'b00101100: delay<=32'h1F240;
	8'b00110101: delay<=32'h1B6A4;
	8'b00111100: delay<=32'h18CB7;
	8'b01000011: delay<=32'h17544;
	8'b01000100: delay<=32'h14C8B;
	8'b01001101: delay<=32'h12843;
	8'b00011110: delay<=32'h2C0A2;
	8'b00100110: delay<=32'h273C2;
	8'b00101110: delay<=32'h20FE1;
	8'b00110110: delay<=32'h1D649;
	8'b00111101: delay<=32'h1A2FA;
	8'b01000110: delay<=32'h16051;
	8'b01000101: delay<=32'h139E1;
	/*
	if(keyboard == 8'b00010101) delay<=32'h2F691;
	else if(keyboard == 8'b00011101) delay<=32'h29AB2;
	else if(keyboard == 8'b00100100) delay<=32'h24A26;
	else if(keyboard == 8'b00101101) delay<=32'h230E4;
	else if(keyboard == 8'b00101100) delay<=32'h1F240;
	else if(keyboard == 8'b00110101) delay<=32'h1B6A4;
	else if(keyboard == 8'b00111100) delay<=32'h18CB7;
	else if(keyboard == 8'b01000011) delay<=32'h17544;
	else if(keyboard == 8'b01000100) delay<=32'h14C8B;
	else if(keyboard == 8'b01001101) delay<=32'h12843;
	else if(keyboard == 8'b00011110) delay<=32'h2C0A2;
	else if(keyboard == 8'b00100110) delay<=32'h273C2;
	else if(keyboard == 8'b00101110) delay<=32'h20FE1;
	else if(keyboard == 8'b00110110) delay<=32'h1D649;
	else if(keyboard == 8'b00111101) delay<=32'h1A2FA;
	else if(keyboard == 8'b01000110) delay<=32'h16051;
	else if(keyboard == 8'b01000101) delay<=32'h139E1;
	else delay<= 32'b1;
	*/
default: delay<=32'b1;
endcase
end
//divinde 50million by each frequerncy


/*****************************************************************************
 *                             Sequential Logic                              *
 *****************************************************************************/

always @(posedge CLOCK_50)
	if(delay_cnt == delay) begin
		delay_cnt <= 0;
		snd <= !snd;
	end else delay_cnt <= delay_cnt + 1;

/*****************************************************************************
 *                            Combinational Logic                            *
 *****************************************************************************/

//assign delay = {SW[3:0], 15'd3000};

wire [31:0] sound = (~(keyboard == 8'b00010101 || keyboard == 8'b00011101 || keyboard == 8'b00100100 || keyboard == 8'b00101101 || keyboard == 8'b00101100 || keyboard == 8'b00110101 || keyboard == 8'b00111100 || keyboard == 8'b01000011 || keyboard == 8'b01000100 || keyboard == 8'b01001101 ||keyboard == 8'b00011110 || keyboard == 8'b00100110 || keyboard == 8'b00101110 || keyboard == 8'b00110110 || keyboard == 8'b00111101 || keyboard == 8'b01000110 || keyboard == 8'b01000101)) ? 0 : snd ? 32'd10000000 : -32'd10000000;


assign read_audio_in			= audio_in_available & audio_out_allowed;

assign left_channel_audio_out	= left_channel_audio_in+sound;
assign right_channel_audio_out	= right_channel_audio_in+sound;
assign write_audio_out			= audio_in_available & audio_out_allowed;

/*****************************************************************************
 *                              Internal Modules                             *
 *****************************************************************************/

Audio_Controller Audio_Controller (
	// Inputs
	.CLOCK_50						(CLOCK_50),
	.reset						(~KEY[0]),

	.clear_audio_in_memory		(),
	.read_audio_in				(read_audio_in),
	
	.clear_audio_out_memory		(),
	.left_channel_audio_out		(left_channel_audio_out),
	.right_channel_audio_out	(right_channel_audio_out),
	.write_audio_out			(write_audio_out),

	.AUD_ADCDAT					(AUD_ADCDAT),

	// Bidirectionals
	.AUD_BCLK					(AUD_BCLK),
	.AUD_ADCLRCK				(AUD_ADCLRCK),
	.AUD_DACLRCK				(AUD_DACLRCK),


	// Outputs
	.audio_in_available			(audio_in_available),
	.left_channel_audio_in		(left_channel_audio_in),
	.right_channel_audio_in		(right_channel_audio_in),

	.audio_out_allowed			(audio_out_allowed),

	.AUD_XCK					(AUD_XCK),
	.AUD_DACDAT					(AUD_DACDAT)

);

avconf #(.USE_MIC_INPUT(1)) avc (
	.FPGA_I2C_SCLK					(FPGA_I2C_SCLK),
	.FPGA_I2C_SDAT					(FPGA_I2C_SDAT),
	.CLOCK_50					(CLOCK_50),
	.reset						(~KEY[0])
);

PS2_Controller c1(
	.CLOCK_50(CLOCK_50),
	.reset(~KEY[0]),

	// Bidirectionals
	.PS2_CLK(PS2_CLK),					// PS2 Clock
 	.PS2_DAT(PS2_DAT),					// PS2 Data

	// Outputs

	.received_data(keyboard),
	.received_data_en(e)
	);
endmodule


